library verilog;
use verilog.vl_types.all;
entity mult_with_3_stages_pipeline_vlg_vec_tst is
end mult_with_3_stages_pipeline_vlg_vec_tst;
